library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SEG_8D is
	PORT(	DATA_A	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DATA_B	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DATA_C	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			DATA_D	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			CLK		: IN STD_LOGIC;
			SEG		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			POS		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
end SEG_8D;

architecture Behavioral of SEG_8D is

	SIGNAL CNT: INTEGER RANGE 0 TO 52083 := 0;
	SIGNAL SHIFT_CLK: STD_LOGIC := '0';
	SIGNAL SHIFT_POS: STD_LOGIC_VECTOR(7 DOWNTO 0) := "11111110";
	SIGNAL VALUE: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	
	COMPONENT BCD is
		PORT(	DATA: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
				SEG: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	end COMPONENT;

begin

	COUNT: PROCESS(CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			CNT <= CNT + 1;
			IF CNT = 52083 THEN
				CNT <= 0;
				SHIFT_CLK <= NOT SHIFT_CLK;
			END IF;
		END IF;
	END PROCESS;
	
	SHIFT: PROCESS(SHIFT_CLK)
	BEGIN
		IF RISING_EDGE(SHIFT_CLK) THEN
			SHIFT_POS <= SHIFT_POS(6 DOWNTO 0) & SHIFT_POS(7);
		END IF;
	END PROCESS;
	
	POS <= SHIFT_POS;
	
	WITH SHIFT_POS SELECT VALUE <=
		DATA_A(7 DOWNTO 4) WHEN "11111110",
		DATA_A(3 DOWNTO 0) WHEN "11111101",
		DATA_B(7 DOWNTO 4) WHEN "11111011",
		DATA_B(3 DOWNTO 0) WHEN "11110111",
		DATA_C(7 DOWNTO 4) WHEN "11101111",
		DATA_C(3 DOWNTO 0) WHEN "11011111",
		DATA_D(7 DOWNTO 4) WHEN "10111111",
		DATA_D(3 DOWNTO 0) WHEN OTHERS;
		
	DIGITS: BCD PORT MAP(
		DATA => VALUE,
		SEG => SEG
	);
	
end Behavioral;

